module delay1(b1,b2);

input wire [1:0] b1;
input wire [1:0] b2;

//register, adder
